module test(
    input   clk,
    input   rst

);

endmodule
