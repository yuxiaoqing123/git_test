module test(
    input   ck,
    input   rst

);

endmodule
